`timescale 1ns / 1ps
/**
	@file GuessGenerator.v
	@author Andrew D. Zonenberg
	@brief Guess generation module
 */
module GuessGenerator(clk, guess);

	input wire clk;
	output reg[63:0] guess;
	

endmodule
